// source_sel_avst_credit_multiplexer_altera_merlin_multiplexer_110_l2uosvi.v

// Generated using ACDS version 21.1 169

`timescale 1 ps / 1 ps
module source_sel_avst_credit_multiplexer_altera_merlin_multiplexer_110_l2uosvi (
		input  wire        clk,                 //       clk.clk
		input  wire        reset,               // clk_reset.reset
		input  wire        src_ready,           //       src.ready
		output wire        src_valid,           //          .valid
		output wire [63:0] src_data,            //          .data
		output wire [1:0]  src_channel,         //          .channel
		output wire        src_startofpacket,   //          .startofpacket
		output wire        src_endofpacket,     //          .endofpacket
		output wire        sink0_ready,         //     sink0.ready
		input  wire        sink0_valid,         //          .valid
		input  wire [1:0]  sink0_channel,       //          .channel
		input  wire [63:0] sink0_data,          //          .data
		input  wire        sink0_startofpacket, //          .startofpacket
		input  wire        sink0_endofpacket,   //          .endofpacket
		output wire        sink1_ready,         //     sink1.ready
		input  wire        sink1_valid,         //          .valid
		input  wire [1:0]  sink1_channel,       //          .channel
		input  wire [63:0] sink1_data,          //          .data
		input  wire        sink1_startofpacket, //          .startofpacket
		input  wire        sink1_endofpacket,   //          .endofpacket
		output wire        sink2_ready,         //     sink2.ready
		input  wire        sink2_valid,         //          .valid
		input  wire [1:0]  sink2_channel,       //          .channel
		input  wire [63:0] sink2_data,          //          .data
		input  wire        sink2_startofpacket, //          .startofpacket
		input  wire        sink2_endofpacket,   //          .endofpacket
		output wire        sink3_ready,         //     sink3.ready
		input  wire        sink3_valid,         //          .valid
		input  wire [1:0]  sink3_channel,       //          .channel
		input  wire [63:0] sink3_data,          //          .data
		input  wire        sink3_startofpacket, //          .startofpacket
		input  wire        sink3_endofpacket    //          .endofpacket
	);

	source_sel_altera_merlin_multiplexer_1921_hjfvwkq mux_inst_name (
		.clk                 (clk),                 //   input,   width = 1,       clk.clk
		.reset               (reset),               //   input,   width = 1, clk_reset.reset
		.src_ready           (src_ready),           //   input,   width = 1,       src.ready
		.src_valid           (src_valid),           //  output,   width = 1,          .valid
		.src_data            (src_data),            //  output,  width = 64,          .data
		.src_channel         (src_channel),         //  output,   width = 2,          .channel
		.src_startofpacket   (src_startofpacket),   //  output,   width = 1,          .startofpacket
		.src_endofpacket     (src_endofpacket),     //  output,   width = 1,          .endofpacket
		.sink0_ready         (sink0_ready),         //  output,   width = 1,     sink0.ready
		.sink0_valid         (sink0_valid),         //   input,   width = 1,          .valid
		.sink0_channel       (sink0_channel),       //   input,   width = 2,          .channel
		.sink0_data          (sink0_data),          //   input,  width = 64,          .data
		.sink0_startofpacket (sink0_startofpacket), //   input,   width = 1,          .startofpacket
		.sink0_endofpacket   (sink0_endofpacket),   //   input,   width = 1,          .endofpacket
		.sink1_ready         (sink1_ready),         //  output,   width = 1,     sink1.ready
		.sink1_valid         (sink1_valid),         //   input,   width = 1,          .valid
		.sink1_channel       (sink1_channel),       //   input,   width = 2,          .channel
		.sink1_data          (sink1_data),          //   input,  width = 64,          .data
		.sink1_startofpacket (sink1_startofpacket), //   input,   width = 1,          .startofpacket
		.sink1_endofpacket   (sink1_endofpacket),   //   input,   width = 1,          .endofpacket
		.sink2_ready         (sink2_ready),         //  output,   width = 1,     sink2.ready
		.sink2_valid         (sink2_valid),         //   input,   width = 1,          .valid
		.sink2_channel       (sink2_channel),       //   input,   width = 2,          .channel
		.sink2_data          (sink2_data),          //   input,  width = 64,          .data
		.sink2_startofpacket (sink2_startofpacket), //   input,   width = 1,          .startofpacket
		.sink2_endofpacket   (sink2_endofpacket),   //   input,   width = 1,          .endofpacket
		.sink3_ready         (sink3_ready),         //  output,   width = 1,     sink3.ready
		.sink3_valid         (sink3_valid),         //   input,   width = 1,          .valid
		.sink3_channel       (sink3_channel),       //   input,   width = 2,          .channel
		.sink3_data          (sink3_data),          //   input,  width = 64,          .data
		.sink3_startofpacket (sink3_startofpacket), //   input,   width = 1,          .startofpacket
		.sink3_endofpacket   (sink3_endofpacket)    //   input,   width = 1,          .endofpacket
	);

endmodule
